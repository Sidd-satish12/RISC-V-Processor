`include "sys_defs.svh"

// -------------------------------------------------------------
// Minimal N-way freelist (mask-driven)
// - Dispatch provides AllocReqMask[N]: which lanes need a tag.
// - Freelist exposes next up to N tags in FreeReg[0..N-1].
//   Dispatch must only consume the first pop_now tags, where
//     pop_now = min(popcount(AllocReqMask), FreeSlotsForN).
// - Retire returns up to N old tags.
// - Optional reseed on mispredict (from Retire) using arch map.
// -------------------------------------------------------------
module freelist #(
    parameter int ALLOC_WIDTH = `N,                // Number of allocation requests per cycle
    parameter int PR_COUNT    = `PHYS_REG_SZ_R10K
) (
    input clock,  // system clock
    input reset,  // system reset

    // From dispatch: allocation requests
    input logic [ALLOC_WIDTH-1:0] alloc_req,  // Request allocation for each dispatch lane

    // From retire: deallocation requests
    input logic [PR_COUNT-1:0] free_mask,  // Bit mask of registers being freed

    // Outputs to dispatch
    output logic [ALLOC_WIDTH-1:0][PR_COUNT-1:0] granted_regs  // Granted physical registers for each allocation request
);

    // Grant matrix from allocator: grants[requester][resource]
    logic [ALLOC_WIDTH-1:0][PR_COUNT-1:0] grants;

    // Allocator instance for physical register allocation
    allocator #(
        .NUM_RESOURCES(PR_COUNT),
        .NUM_REQUESTS (ALLOC_WIDTH)
    ) reg_allocator (
        .reset(reset),
        .clock(clock),
        .req  (alloc_req),  // Allocation requests
        .clear(free_mask),  // Registers being freed
        .grant(grants)      // Grant matrix
    );

    // Output grant matrix directly
    assign granted_regs = grants;

endmodule
