`include "sys_defs.svh"

// Basic testbench for stage_issue module
// Tests basic functionality for synthesis verification

module testbench;

    logic clock, reset;
    logic mispredict;
    logic failed;

    // Inputs to stage_issue
    RS_BANKS rs_banks;
    FU_GRANTS fu_grants;

    // Outputs from stage_issue
    ISSUE_CLEAR issue_clear;
    ISSUE_ENTRIES issue_entries;

    stage_issue dut (
        .clock(clock),
        .reset(reset),
        .mispredict(mispredict),
        .rs_banks(rs_banks),
        .fu_grants(fu_grants),
        .issue_clear(issue_clear),
        .issue_entries(issue_entries)
    );

    always begin
        #50 clock = ~clock;  // 100ns period
    end

    // Helper function to create a default empty entry
    function RS_ENTRY empty_entry;
        empty_entry.valid = 0;
        empty_entry.opa_select = OPA_IS_RS1;
        empty_entry.opb_select = OPB_IS_RS2;
        empty_entry.op_type = OP_ALU_ADD;
        empty_entry.src1_tag = 0;
        empty_entry.src1_ready = 0;
        empty_entry.src1_value = 0;
        empty_entry.src2_tag = 0;
        empty_entry.src2_ready = 0;
        empty_entry.src2_value = 0;
        empty_entry.dest_tag = 0;
        empty_entry.rob_idx = 0;
        empty_entry.rob_wrap = 0;
        empty_entry.PC = 0;
        empty_entry.pred_taken = 0;
        empty_entry.pred_target = 0;
    endfunction

    // Helper function to create a ready ALU entry
    function RS_ENTRY ready_alu_entry(input int rob_idx_val, input int rob_wrap_val = 0);
        ready_alu_entry = empty_entry();
        ready_alu_entry.valid = 1;
        ready_alu_entry.op_type.category = CAT_ALU;
        ready_alu_entry.op_type.func = ADD;
        ready_alu_entry.src1_ready = 1;
        ready_alu_entry.src2_ready = 1;
        ready_alu_entry.rob_idx = rob_idx_val;
        ready_alu_entry.rob_wrap = rob_wrap_val;
    endfunction

    // Helper function to create a ready MULT entry
    function RS_ENTRY ready_mult_entry(input int rob_idx_val, input int rob_wrap_val = 0);
        ready_mult_entry = empty_entry();
        ready_mult_entry.valid = 1;
        ready_mult_entry.op_type.category = CAT_MULT;
        ready_mult_entry.op_type.func = MUL;
        ready_mult_entry.src1_ready = 1;
        ready_mult_entry.src2_ready = 1;
        ready_mult_entry.rob_idx = rob_idx_val;
        ready_mult_entry.rob_wrap = rob_wrap_val;
    endfunction

    // Helper function to create a ready BRANCH entry
    function RS_ENTRY ready_branch_entry(input int rob_idx_val, input int rob_wrap_val = 0);
        ready_branch_entry = empty_entry();
        ready_branch_entry.valid = 1;
        ready_branch_entry.op_type.category = CAT_BRANCH;
        ready_branch_entry.op_type.func = EQ;
        ready_branch_entry.src1_ready = 1;
        ready_branch_entry.src2_ready = 1;
        ready_branch_entry.rob_idx = rob_idx_val;
        ready_branch_entry.rob_wrap = rob_wrap_val;
    endfunction

    // Helper function to create a ready MEM entry
    function RS_ENTRY ready_mem_entry(input int rob_idx_val, input int rob_wrap_val = 0);
        ready_mem_entry = empty_entry();
        ready_mem_entry.valid = 1;
        ready_mem_entry.op_type.category = CAT_MEM;
        ready_mem_entry.op_type.func = LOAD_WORD;
        ready_mem_entry.src1_ready = 1;
        ready_mem_entry.src2_ready = 1;
        ready_mem_entry.rob_idx = rob_idx_val;
        ready_mem_entry.rob_wrap = rob_wrap_val;
    endfunction

    // Helper function to create a not-ready entry
    function RS_ENTRY not_ready_entry(input OP_CATEGORY cat, input int rob_idx_val);
        not_ready_entry = empty_entry();
        not_ready_entry.valid = 1;
        not_ready_entry.op_type.category = cat;
        not_ready_entry.src1_ready = 0;
        not_ready_entry.src2_ready = 0;
        not_ready_entry.rob_idx = rob_idx_val;
    endfunction

    // Helper to print issue results
    task print_issue_results(input string label);
        $display("\n=== %s ===", label);
        $display("ALU clears: valid=%b, idxs=%p", issue_clear.valid_alu, issue_clear.idxs_alu);
        $display("MULT clears: valid=%b, idxs=%p", issue_clear.valid_mult, issue_clear.idxs_mult);
        $display("BRANCH clears: valid=%b, idxs=%p", issue_clear.valid_branch, issue_clear.idxs_branch);
        $display("MEM clears: valid=%b, idxs=%p", issue_clear.valid_mem, issue_clear.idxs_mem);
        $display("");
    endtask

    // Helper to reset and wait for proper timing
    task reset_dut;
        reset = 1;
        @(negedge clock);
        @(negedge clock);
        reset = 0;
        @(negedge clock);
    endtask

    initial begin
        int test_num = 1;
        clock = 0;
        reset = 1;
        failed = 0;
        mispredict = 0;

        // Initialize inputs
        rs_banks = '0;
        fu_grants = '0;

        reset_dut();

        // Test 1: Single ready ALU instruction, FU available
        $display("\nTest %0d: Single ready ALU instruction, FU available", test_num++);
        reset_dut();
        begin
            logic any_alu_clear;
            rs_banks = '0;
            rs_banks.alu[0] = ready_alu_entry(10);
            fu_grants = '0;
            fu_grants.alu = {`NUM_FU_ALU{1'b1}};

            // Wait for allocator to stabilize (may need a cycle)
            @(posedge clock);
            #10;
            @(posedge clock);
            #10;

            // Check that an ALU entry was issued
            any_alu_clear = |issue_clear.valid_alu;
            if (any_alu_clear) begin
                $display("  PASS: ALU clear valid is set");
            end else begin
                $display("  FAIL: ALU clear valid should be set");
                failed = 1;
            end
        end

        // Test 2: Single ready MULT instruction, FU available
        $display("\nTest %0d: Single ready MULT instruction, FU available", test_num++);
        reset_dut();
        begin
            logic any_mult_clear;
            rs_banks = '0;
            rs_banks.mult[0] = ready_mult_entry(15);
            fu_grants = '0;
            fu_grants.mult = {`NUM_FU_MULT{1'b1}};

            @(posedge clock);
            #10;
            @(posedge clock);
            #10;

            any_mult_clear = |issue_clear.valid_mult;
            if (any_mult_clear) begin
                $display("  PASS: MULT clear valid is set");
            end else begin
                $display("  FAIL: MULT clear valid should be set");
                failed = 1;
            end
        end

        // Test 3: Single ready BRANCH instruction, FU available
        $display("\nTest %0d: Single ready BRANCH instruction, FU available", test_num++);
        reset_dut();
        begin
            logic any_branch_clear;
            rs_banks = '0;
            rs_banks.branch[0] = ready_branch_entry(20);
            fu_grants = '0;
            fu_grants.branch = {`NUM_FU_BRANCH{1'b1}};

            @(posedge clock);
            #10;
            @(posedge clock);
            #10;

            any_branch_clear = |issue_clear.valid_branch;
            if (any_branch_clear) begin
                $display("  PASS: BRANCH clear valid is set");
            end else begin
                $display("  FAIL: BRANCH clear valid should be set");
                failed = 1;
            end
        end

        // Test 4: Single ready MEM instruction, FU available
        $display("\nTest %0d: Single ready MEM instruction, FU available", test_num++);
        reset_dut();
        begin
            logic any_mem_clear;
            rs_banks = '0;
            rs_banks.mem[0] = ready_mem_entry(25);
            fu_grants = '0;
            fu_grants.mem = {`NUM_FU_MEM{1'b1}};

            @(posedge clock);
            #10;
            @(posedge clock);
            #10;

            any_mem_clear = |issue_clear.valid_mem;
            if (any_mem_clear) begin
                $display("  PASS: MEM clear valid is set");
            end else begin
                $display("  FAIL: MEM clear valid should be set");
                failed = 1;
            end
        end

        // Test 5: Multiple ready instructions across categories
        $display("\nTest %0d: Multiple ready instructions across categories", test_num++);
        reset_dut();
        begin
            logic any_alu, any_mult, any_branch, any_mem;
            rs_banks = '0;
            rs_banks.alu[0] = ready_alu_entry(10);
            rs_banks.mult[0] = ready_mult_entry(15);
            rs_banks.branch[0] = ready_branch_entry(20);
            rs_banks.mem[0] = ready_mem_entry(25);
            fu_grants = '0;
            fu_grants.alu = {`NUM_FU_ALU{1'b1}};
            fu_grants.mult = {`NUM_FU_MULT{1'b1}};
            fu_grants.branch = {`NUM_FU_BRANCH{1'b1}};
            fu_grants.mem = {`NUM_FU_MEM{1'b1}};

            @(posedge clock);
            #10;
            @(posedge clock);
            #10;

            // Check that all categories issued
            any_alu = |issue_clear.valid_alu;
            any_mult = |issue_clear.valid_mult;
            any_branch = |issue_clear.valid_branch;
            any_mem = |issue_clear.valid_mem;
            if (any_alu && any_mult && any_branch && any_mem) begin
                $display("  PASS: All categories issued");
            end else begin
                $display("  FAIL: All categories should issue (alu=%b, mult=%b, branch=%b, mem=%b)", any_alu, any_mult,
                         any_branch, any_mem);
                failed = 1;
            end
        end

        // Test 6: Not-ready instruction should not issue
        $display("\nTest %0d: Not-ready instruction should not issue", test_num++);
        reset_dut();
        begin
            logic any_alu_clear;
            rs_banks = '0;
            rs_banks.alu[0] = not_ready_entry(CAT_ALU, 10);
            fu_grants = '0;
            fu_grants.alu = {`NUM_FU_ALU{1'b1}};

            @(posedge clock);
            #10;
            @(posedge clock);
            #10;

            any_alu_clear = |issue_clear.valid_alu;
            if (!any_alu_clear) begin
                $display("  PASS: Not-ready instruction did not issue");
            end else begin
                $display("  FAIL: Not-ready instruction should not issue");
                failed = 1;
            end
        end

        // Test 7: Invalid entry should not issue
        $display("\nTest %0d: Invalid entry should not issue", test_num++);
        reset_dut();
        begin
            logic any_alu_clear;
            rs_banks = '0;
            rs_banks.alu[0] = empty_entry();  // Invalid
            fu_grants = '0;
            fu_grants.alu = {`NUM_FU_ALU{1'b1}};

            @(posedge clock);
            #10;
            @(posedge clock);
            #10;

            any_alu_clear = |issue_clear.valid_alu;
            if (!any_alu_clear) begin
                $display("  PASS: Invalid entry did not issue");
            end else begin
                $display("  FAIL: Invalid entry should not issue");
                failed = 1;
            end
        end

        // Test 8: No FU available should not issue
        $display("\nTest %0d: No FU available should not issue", test_num++);
        reset_dut();
        begin
            logic any_alu_clear;
            rs_banks = '0;
            rs_banks.alu[0] = ready_alu_entry(10);
            fu_grants = '0;
            fu_grants.alu = {`NUM_FU_ALU{1'b0}};  // No FUs available

            @(posedge clock);
            #10;
            @(posedge clock);
            #10;

            any_alu_clear = |issue_clear.valid_alu;
            if (!any_alu_clear) begin
                $display("  PASS: No issue when no FU available");
            end else begin
                $display("  FAIL: Should not issue when no FU available");
                failed = 1;
            end
        end

        // Test 9: Reset clears issue register
        $display("\nTest %0d: Reset clears issue register", test_num++);
        reset_dut();
        begin
            rs_banks = '0;
            rs_banks.alu[0] = ready_alu_entry(10);
            fu_grants = '0;
            fu_grants.alu = {`NUM_FU_ALU{1'b1}};

            @(posedge clock);
            #10;

            // Apply reset
            reset = 1;
            @(posedge clock);
            #10;

            // Check that issue register is cleared
            if (issue_entries.alu[0].valid == 0) begin
                $display("  PASS: Reset clears issue register");
            end else begin
                $display("  FAIL: Reset should clear issue register");
                failed = 1;
            end
        end

        // Test 10: Mispredict clears issue register
        $display("\nTest %0d: Mispredict clears issue register", test_num++);
        reset_dut();
        begin
            rs_banks = '0;
            rs_banks.alu[0] = ready_alu_entry(10);
            fu_grants = '0;
            fu_grants.alu = {`NUM_FU_ALU{1'b1}};

            @(posedge clock);
            #10;

            // Apply mispredict
            mispredict = 1;
            @(posedge clock);
            #10;

            // Check that issue register is cleared
            if (issue_entries.alu[0].valid == 0) begin
                $display("  PASS: Mispredict clears issue register");
            end else begin
                $display("  FAIL: Mispredict should clear issue register");
                failed = 1;
            end
        end

        // Test 11: Multiple ALU instructions, multiple FUs
        $display("\nTest %0d: Multiple ALU instructions, multiple FUs", test_num++);
        reset_dut();
        begin
            int count;
            int i;
            rs_banks = '0;
            rs_banks.alu[0] = ready_alu_entry(10);
            rs_banks.alu[1] = ready_alu_entry(15);
            rs_banks.alu[2] = ready_alu_entry(20);
            fu_grants = '0;
            fu_grants.alu = {`NUM_FU_ALU{1'b1}};

            @(posedge clock);
            #10;
            @(posedge clock);
            #10;

            // Check that multiple entries can be issued
            count = 0;
            for (i = 0; i < `NUM_FU_ALU; i++) begin
                if (issue_clear.valid_alu[i]) count++;
            end
            if (count > 0 && count <= `NUM_FU_ALU) begin
                $display("  PASS: Issued %0d ALU instructions", count);
            end else begin
                $display("  FAIL: Should issue between 1 and %0d ALU instructions, got %0d", `NUM_FU_ALU, count);
                failed = 1;
            end
        end

        $display("\n");
        if (failed) begin
            $display("@@@ FAILED");
        end else begin
            $display("@@@ PASSED");
        end

        $finish;
    end

endmodule
