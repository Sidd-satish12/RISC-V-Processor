/////////////////////////////////////////////////////////////////////////
//                                                                     //
//   Modulename :  cpu_test.sv                                         //
//                                                                     //
//  Description :  Testbench module for the VeriSimpleV processor.     //
//                                                                     //
/////////////////////////////////////////////////////////////////////////

`include "sys_defs.svh"

// P4 TODO: Add your own debugging framework. Basic printing of data structures
//          is an absolute necessity for the project. You can use C functions 
//          like in test/pipeline_print.c or just do everything in verilog.
//          Be careful about running out of space on CAEN printing lots of state
//          for longer programs (alexnet, outer_product, etc.)

// These link to the pipeline_print.c file in this directory, and are used below to print
// detailed output to the pipeline_output_file, initialized by open_pipeline_output_file()
import "DPI-C" function string decode_inst(int inst);
// Pipeline printing disabled for OOO processor
// import "DPI-C" function void open_pipeline_output_file(string file_name);
// import "DPI-C" function void print_header();
// import "DPI-C" function void print_cycles(int clock_count);
// import "DPI-C" function void print_stage(
//     int inst,
//     int npc,
//     int valid_inst
// );
// import "DPI-C" function void print_reg(
//     int wb_data,
//     int wb_idx,
//     int wb_en
// );
// import "DPI-C" function void print_membus(int proc2mem_command, int proc2mem_addr,
//                                           int proc2mem_data_hi, int proc2mem_data_lo);
// import "DPI-C" function void close_pipeline_output_file();


`define TB_MAX_CYCLES 20


module testbench;
    // string inputs for loading memory and output files
    // run like: cd build && ./simv +MEMORY=../programs/mem/<my_program>.mem +OUTPUT=../output/<my_program>
    // this testbench will generate 4 output files based on the output
    // named OUTPUT.{out cpi, wb, ppln} for the memory, cpi, writeback, and pipeline outputs.
    string program_memory_file, output_name;
    string out_outfile, cpi_outfile, writeback_outfile;  //, pipeline_outfile;
    int out_fileno, cpi_fileno, wb_fileno;  // verilog uses integer file handles with $fopen and $fclose

    // variables used in the testbench
    logic                                 clock;
    logic                                 reset;
    logic              [            31:0] clock_count;  // also used for terminating infinite loops
    logic              [            31:0] instr_count;

    // Disconnected: proc2mem/mem2proc portions (fake-fetch)
    // MEM_COMMAND             proc2mem_command;
    // ADDR                    proc2mem_addr;
    // MEM_BLOCK               proc2mem_data;
    // MEM_TAG                 mem2proc_transaction_tag;
    // MEM_BLOCK               mem2proc_data;
    // MEM_TAG                 mem2proc_data_tag;
    // MEM_SIZE                proc2mem_size;

    COMMIT_PACKET      [          `N-1:0] committed_insts;
    EXCEPTION_CODE                        error_status = NO_ERROR;

    ADDR                                  if_NPC_dbg;
    DATA                                  if_inst_dbg;
    logic                                 if_valid_dbg;
    ADDR                                  if_id_NPC_dbg;
    DATA                                  if_id_inst_dbg;
    logic                                 if_id_valid_dbg;
    ADDR                                  id_ex_NPC_dbg;
    DATA                                  id_ex_inst_dbg;
    logic                                 id_ex_valid_dbg;
    ADDR                                  ex_mem_NPC_dbg;
    DATA                                  ex_mem_inst_dbg;
    logic                                 ex_mem_valid_dbg;
    ADDR                                  mem_wb_NPC_dbg;
    DATA                                  mem_wb_inst_dbg;
    logic                                 mem_wb_valid_dbg;

    // OOO debug signals
    logic              [          `N-1:0] rob_head_valids;
    ROB_ENTRY          [          `N-1:0] rob_head_entries;
    logic              [$clog2(`N+1)-1:0] dispatch_count;
    RS_GRANTED_BANKS                      rs_granted;

    // Additional debug for RS and issue state
    logic              [  `RS_ALU_SZ-1:0] rs_alu_ready;
    ISSUE_ENTRIES                         issue_entries;

    // Execute stage debug signals
    logic              [          `N-1:0] ex_valid;
    EX_COMPLETE_PACKET                    ex_comp;

    // Complete stage debug signals
    ROB_UPDATE_PACKET                     rob_update_packet;

    // ----------------------------------------------------------------
    // Fake-Fetch wires (testbench <-> cpu)
    // ----------------------------------------------------------------
    ADDR                                  fake_pc;
    DATA                                  fake_instr                                               [`N-1:0];
    logic              [$clog2(`N+1)-1:0] fake_nvalid;
    logic              [$clog2(`N+1)-1:0] fake_consumed;

    logic                                 ff_branch_taken;
    ADDR                                  ff_branch_target;

    // Debug Output PRF
    DATA [`PHYS_REG_SZ_R10K-1:0] regfile_entries;

    // Debug output Architecture map table
    MAP_ENTRY [`ARCH_REG_SZ-1:0] arch_table_snapshot;

    // debug output rs_alu
    RS_ENTRY            [   `RS_ALU_SZ-1:0] rs_alu_entries;


    // Instantiate the Pipeline
    cpu verisimpleV (
        // Inputs
        .clock(clock),
        .reset(reset),
        // Disconnected: mem2proc portions (fake-fetch)
        // .mem2proc_transaction_tag(mem2proc_transaction_tag),
        // .mem2proc_data           (mem2proc_data),
        // .mem2proc_data_tag       (mem2proc_data_tag),

        // Disconnected: proc2mem portions (fake-fetch)
        // .proc2mem_command(proc2mem_command),
        // .proc2mem_addr   (proc2mem_addr),
        // .proc2mem_data   (proc2mem_data),
        // `ifndef CACHE_MODE
        // .proc2mem_size   (proc2mem_size),
        // `endif

        .committed_insts(committed_insts),

        .fetch_NPC_dbg     (if_NPC_dbg),
        .fetch_inst_dbg    (if_inst_dbg),
        .fetch_valid_dbg   (if_valid_dbg),
        .dispatch_NPC_dbg  (if_id_NPC_dbg),
        .dispatch_inst_dbg (if_id_inst_dbg),
        .dispatch_valid_dbg(if_id_valid_dbg),
        .issue_NPC_dbg     (id_ex_NPC_dbg),
        .issue_inst_dbg    (id_ex_inst_dbg),
        .issue_valid_dbg   (id_ex_valid_dbg),
        .execute_NPC_dbg   (ex_mem_NPC_dbg),
        .execute_inst_dbg  (ex_mem_inst_dbg),
        .execute_valid_dbg (ex_mem_valid_dbg),
        .complete_NPC_dbg  (mem_wb_NPC_dbg),    // Using old names for compatibility
        .complete_inst_dbg (mem_wb_inst_dbg),
        .complete_valid_dbg(mem_wb_valid_dbg),
        .retire_NPC_dbg    (),                  // Not used in testbench
        .retire_inst_dbg   (),
        .retire_valid_dbg  (),

        // Additional debug outputs
        .rob_head_valids_dbg(rob_head_valids),
        .rob_head_entries_dbg(rob_head_entries),
        .dispatch_count_dbg(dispatch_count),
        .rs_granted_dbg(rs_granted),
        .rs_alu_ready_dbg(rs_alu_ready),
        .issue_entries_dbg(issue_entries),

        // Execute stage debug outputs
        .ex_valid_dbg(ex_valid),
        .ex_comp_dbg (ex_comp),

        // Complete stage debug outputs
        .rob_update_packet_dbg(rob_update_packet),

        // Debug output from PRF
        .regfile_entries(regfile_entries),

        // Debug output from architecture map table
        .arch_table_snapshot(arch_table_snapshot),

        // Debug output from RS_ALU
        .rs_alu_entries(rs_alu_entries),

        // ---- Fake-Fetch interface ----
        .ff_instr       (fake_instr),
        .ff_pc          (fake_pc),
        .ff_nvalid      (fake_nvalid),
        .ff_consumed    (fake_consumed),
        .branch_taken_o (ff_branch_taken),
        .branch_target_o(ff_branch_target)
    );


    // Instruction Memory (for fake-fetch only - data operations disconnected)
    mem memory (
        // Only connect clock for initialization
        .clock           (clock),
        // Data operations disconnected
        .proc2mem_command(MEM_NONE),
        .proc2mem_addr   ('0),
        .proc2mem_data   ('0),
`ifndef CACHE_MODE
        .proc2mem_size   (DOUBLE),
`endif

        // Outputs not used for fake-fetch
        .mem2proc_transaction_tag(),
        .mem2proc_data           (),
        .mem2proc_data_tag       ()
    );


    // Generate System Clock
    always begin
        #(`CLOCK_PERIOD / 2.0);
        clock = ~clock;
    end

    // ----------------------------------------------------------------
    // Fake-Fetch: PC register
    // ----------------------------------------------------------------
    always_ff @(posedge clock) begin
        if (reset) begin
            fake_pc <= '0;
        end else begin
            if (ff_branch_taken) begin
                fake_pc <= ff_branch_target;
            end else begin
                // Advance by 4*X where X = fake_consumed from CPU
                fake_pc <= fake_pc + 32'(4 * fake_consumed);
            end
        end
    end

    // ----------------------------------------------------------------
    // Read a 32b instruction from unified memory at byte address 'addr'
    // ----------------------------------------------------------------
    function DATA get_inst32(input ADDR addr);
        MEM_BLOCK blk;
        begin
            blk = memory.unified_memory[addr[31:3]];  // 8B-aligned line
            get_inst32 = blk.word_level[addr[2]];  // 0: low word, 1: high word
        end
    endfunction

    // ----------------------------------------------------------------
    // Build the N-wide bundle every cycle (sequential @ fake_pc + 4*i)
    // ----------------------------------------------------------------
    int count;
    always_comb begin
        count = 0;
        for (int i = 0; i < `N; i++) begin
            fake_instr[i] = get_inst32(fake_pc + 32'(4 * i));
            if (fake_instr[i] != 32'b0) begin
                count++;
            end
        end
        fake_nvalid = count;  // simple model: always provide N; CPU decides how many to take
    end


    initial begin
        $dumpfile("cpu_test.vcd");
        $dumpvars(0, testbench);

        $display("\n---- Starting CPU Testbench (Fake-Fetch) ----\n");

        // set paramterized strings, see comment at start of module
        if ($value$plusargs("MEMORY=%s", program_memory_file)) begin
            $display("Using memory file  : %s", program_memory_file);
        end else begin
            $display("Did not receive '+MEMORY=' argument. Exiting.\n");
            $finish;
        end
        if ($value$plusargs("OUTPUT=%s", output_name)) begin
            $display("Using output files : %s.{out, cpi, wb}", output_name);
            out_outfile       = {output_name, ".out"};  // this is how you concatenate strings in verilog
            cpi_outfile       = {output_name, ".cpi"};
            writeback_outfile = {output_name, ".wb"};
            // pipeline_outfile  = {output_name, ".ppln"};
        end else begin
            $display("\nDid not receive '+OUTPUT=' argument. Exiting.\n");
            $finish;
        end

        clock = 1'b0;
        reset = 1'b0;

        $display("\n  %16t : Asserting Reset", $realtime);
        reset = 1'b1;

        @(posedge clock);
        @(posedge clock);

        $display("  %16t : Loading Unified Memory", $realtime);
        // load the compiled program's hex data into the memory module
        $readmemh(program_memory_file, memory.unified_memory);

        @(posedge clock);
        @(posedge clock);
        #1;  // This reset is at an odd time to avoid the pos & neg clock edges
        $display("  %16t : Deasserting Reset", $realtime);
        reset = 1'b0;

        wb_fileno = $fopen(writeback_outfile);
        $fdisplay(wb_fileno, "Register writeback output (hexadecimal)");

        // Pipeline output disabled for OOO processor
        // open_pipeline_output_file(pipeline_outfile);
        // print_header();

        out_fileno = $fopen(out_outfile);

        $display("  %16t : Running Processor", $realtime);
    end


    always @(negedge clock) begin
        if (reset) begin
            // Count the number of cycles and number of instructions committed
            clock_count = 0;
            instr_count = 0;
        end else begin
            #2;  // wait a short time to avoid a clock edge


            clock_count = clock_count + 1;

            if ((clock_count % 10000) == 0) $display("  %16t : %0d cycles", $realtime, clock_count);

            // Optional: peek at fake-fetch behavior
            $display("%0t [FF] pc=%h consumed=%0d br=%0d tgt=%h", $time, fake_pc, fake_consumed, ff_branch_taken,
                     ff_branch_target);

            // Pipeline printing disabled for OOO processor
            // print_cycles(clock_count - 1);
            // print_stage(if_inst_dbg, if_NPC_dbg, {31'b0, if_valid_dbg});  // Fetch
            // print_stage(if_id_inst_dbg, if_id_NPC_dbg, {31'b0, if_id_valid_dbg});  // Dispatch
            // print_stage(id_ex_inst_dbg, id_ex_NPC_dbg, {31'b0, id_ex_valid_dbg});  // Issue
            // print_stage(ex_mem_inst_dbg, ex_mem_NPC_dbg, {31'b0, ex_mem_valid_dbg});  // Execute
            // print_stage(mem_wb_inst_dbg, mem_wb_NPC_dbg, {31'b0, mem_wb_valid_dbg});  // Complete/Retire
            // print_reg(committed_insts[0].data, {27'b0, committed_insts[0].reg_idx}, {31'b0, committed_insts[0].valid});
            // print_membus({30'b0,proc2mem_command}, proc2mem_addr[31:0],
            //              proc2mem_data[63:32], proc2mem_data[31:0]);

            print_custom_data();

            output_reg_writeback_and_maybe_halt();

           
            // Optional: print CDB broadcasts
            for (int i = 0; i < `N; i++) begin
                $display("  CDB[%0d]: valid=%b, tag=%0d, data=%h", i, verisimpleV.cdb_output[i].valid, verisimpleV.cdb_output[i].tag, verisimpleV.cdb_output[i].data);
            end


            // stop the processor
            if (error_status != NO_ERROR || clock_count > `TB_MAX_CYCLES) begin

                $display("  %16t : Processor Finished", $realtime);

                // close the writeback output file (pipeline output disabled)
                // close_pipeline_output_file();
                $fclose(wb_fileno);

                // display the final memory and status
                show_final_mem_and_status(error_status);
                // output the final CPI
                output_cpi_file();

                $display("\n---- Finished CPU Testbench (Fake-Fetch) ----\n");

                #100 $finish;
            end
        end  // if(reset)
    end


    // Task to output register writeback data and potentially halt the processor.
    task output_reg_writeback_and_maybe_halt;
        ADDR pc;
        DATA inst;
        MEM_BLOCK block;
        for (int n = 0; n < `N; n++) begin
            if (committed_insts[n].valid) begin
                // update the count for every committed instruction
                instr_count = instr_count + 1;

                pc = committed_insts[n].NPC - 4;
                block = memory.unified_memory[pc[31:3]];
                inst = block.word_level[pc[2]];
                // print the committed instructions to the writeback output file
                if (committed_insts[n].reg_idx == `ZERO_REG) begin
                    $fdisplay(wb_fileno, "PC %4x:%-8s| ---", pc, decode_inst(inst));
                end else begin
                    $fdisplay(wb_fileno, "PC %4x:%-8s| r%02d=%-8x", pc, decode_inst(inst), committed_insts[n].reg_idx,
                              committed_insts[n].data);
                end

                // exit if we have an illegal instruction or a halt
                if (committed_insts[n].illegal) begin
                    error_status = ILLEGAL_INST;
                    break;
                end else if (committed_insts[n].halt) begin
                    error_status = HALTED_ON_WFI;
                    break;
                end
            end  // if valid
        end
    endtask  // task output_reg_writeback_and_maybe_halt


    // Task to output the final CPI and # of elapsed clock edges
    task output_cpi_file;
        real cpi;
        begin
            cpi = $itor(clock_count) / instr_count;  // must convert int to real
            cpi_fileno = $fopen(cpi_outfile);
            $fdisplay(cpi_fileno, "@@@  %0d cycles / %0d instrs = %f CPI", clock_count, instr_count, cpi);
            $fdisplay(cpi_fileno, "@@@  %4.2f ns total time to execute", clock_count * `CLOCK_PERIOD);
            $fclose(cpi_fileno);
        end
    endtask  // task output_cpi_file


    // Show contents of Unified Memory in both hex and decimal
    // Also output the final processor status
    task show_final_mem_and_status;
        input EXCEPTION_CODE final_status;
        int showing_data;
        begin
            $fdisplay(out_fileno, "\nFinal memory state and exit status:\n");
            $fdisplay(out_fileno, "@@@ Unified Memory contents hex on left, decimal on right: ");
            $fdisplay(out_fileno, "@@@");
            showing_data = 0;
            for (int k = 0; k <= `MEM_64BIT_LINES - 1; k = k + 1) begin
                if (memory.unified_memory[k] != 0) begin
                    $fdisplay(out_fileno, "@@@ mem[%5d] = %x : %0d", k * 8, memory.unified_memory[k], memory.unified_memory[k]);
                    showing_data = 1;
                end else if (showing_data != 0) begin
                    $fdisplay(out_fileno, "@@@");
                    showing_data = 0;
                end
            end
            $fdisplay(out_fileno, "@@@");

            case (final_status)
                LOAD_ACCESS_FAULT: $fdisplay(out_fileno, "@@@ System halted on memory error");
                HALTED_ON_WFI:     $fdisplay(out_fileno, "@@@ System halted on WFI instruction");
                ILLEGAL_INST:      $fdisplay(out_fileno, "@@@ System halted on illegal instruction");
                default:           $fdisplay(out_fileno, "@@@ System halted on unknown error code %x", final_status);
            endcase
            $fdisplay(out_fileno, "@@@");
            $fclose(out_fileno);
        end
    endtask  // task show_final_mem_and_status



    // OPTIONAL: Print our your data here
    // It will go to the $program.log file
    // task print_custom_data;
    //     $display(
    //         "%3d: ROB head valid=%b | Dispatch count=%0d | RS ready=%b | Issue ALU valid=%b | Execute valid=%b | ROB update valid=%b | Committed halt=%b valid=%b",
    //         clock_count - 1, rob_head_valids, dispatch_count, rs_alu_ready, issue_entries.alu[0].valid, ex_valid,
    //         rob_update_packet.valid, committed_insts[0].halt, committed_insts[0].valid);
    // endtask

    task print_custom_data;
        $display("\n--- Cycle %0d ---", clock_count-1);
        $display("ROB head valid: %b | Dispatch count: %0d | RS ALU ready: %b",
                rob_head_valids, dispatch_count, rs_alu_ready);
        
        // Print all ALU RS entries
        // for (int i = 0; i < `RS_ALU_SZ; i++) begin
        //     $display("RS[%0d]: valid=%b ready=%b opcode=%h dest_pr=%0d src_tags=%0d,%0d",
        //             i,
        //             verisimpleV.rs_alu[i].valid,
        //             verisimpleV.rs_alu[i].ready,
        //             verisimpleV.rs_alu[i].opcode,
        //             verisimpleV.rs_alu[i].dest_pr,
        //             verisimpleV.rs_alu[i].src_tag1,
        //             verisimpleV.rs_alu[i].src_tag2);
        // end

        // Print which RS entries were granted to issue
        for (int i = 0; i < `N; i++) begin
            $display("RS grant[%0d]: granted=%b", i, rs_granted.alu[i]);
        end

        // Print Issue entries
        for (int i = 0; i < `N; i++) begin
            $display("Issue entry[%0d]: valid=%b", i, issue_entries.alu[i].valid);
        end

        // Print execution stage
        for (int i = 0; i < `N; i++) begin
            $display("EX[%0d]: valid=%b", i, ex_valid[i]);
        end

        // Print ROB head entries
        for (int i = 0; i < `N; i++) begin
            $display("ROB[%0d]: valid=%b", i, rob_head_valids[i]);
        end

        // Optional: print CDB broadcasts
        for (int i = 0; i < `N; i++) begin
            $display("CDB[%0d]: valid=%b tag=%0d data=%h",
                    i,
                    verisimpleV.cdb_output[i].valid,
                    verisimpleV.cdb_output[i].tag,
                    verisimpleV.cdb_output[i].data);
        end

        for (int i = 0; i < `N; i++) begin
            if (committed_insts[i].valid) begin
                //ADDR pc = committed_insts[i].NPC - 4;
                //string inst_str = decode_inst(get_inst32(pc));
                if (committed_insts[i].reg_idx == `ZERO_REG)
                    $display("COMMIT[%0d]: PC=%h | ---", i, committed_insts[i].NPC - 4);
                else
                    $display("COMMIT[%0d]: PC=%h | r%0d=%h",
                            i, committed_insts[i].NPC - 4, committed_insts[i].reg_idx, committed_insts[i].data);
            end
        end

        //$display("PRF REGISTER 1: %d", regfile_entries[arch_table_snapshot[1].phys_reg]);
        //$display("ARCH MAP TABLE R1 MAPPING ->: %d",arch_table_snapshot[1].phys_reg);

        for (int i = 0; i < `RS_ALU_SZ; i++) begin
            $display("RS[%0d]: valid=%b, opa=%0d, opb=%0d, op_type=%0d, src1_tag=%0d, src1_ready=%b, src2_tag=%0d, src2_ready=%b, dest_tag=%0d, rob_idx=%0d, PC=0x%08h",
                    i,
                    rs_alu_entries[i].valid,
                    rs_alu_entries[i].opa_select,
                    rs_alu_entries[i].opb_select,
                    rs_alu_entries[i].op_type,
                    rs_alu_entries[i].src1_tag,
                    rs_alu_entries[i].src1_ready,
                    rs_alu_entries[i].src2_tag,
                    rs_alu_entries[i].src2_ready,
                    rs_alu_entries[i].dest_tag,
                    rs_alu_entries[i].rob_idx,
                    rs_alu_entries[i].PC
            );
        end

    endtask


endmodule  // module testbench
