module LFSR #(
    parameter NUM_BITS
) (
    input clock,
    input reset,

    input  [NUM_BITS-1:0] seed_data,
    output [NUM_BITS-1:0] data_out
);

    logic [NUM_BITS-1:0] LFSR;
    logic                r_XNOR;

    always @(posedge clock) begin
        if (reset) LFSR <= seed_data;
        else LFSR <= {LFSR[NUM_BITS-1:1], r_XNOR};
    end

    always @(*) begin
        case (NUM_BITS)
            3: begin
                r_XNOR = LFSR[3] ^~ LFSR[2];
            end
            4: begin
                r_XNOR = LFSR[4] ^~ LFSR[3];
            end
            5: begin
                r_XNOR = LFSR[5] ^~ LFSR[3];
            end
            // 6: begin
            //     r_XNOR = LFSR[6] ^~ LFSR[5];
            // end
            // 7: begin
            //     r_XNOR = LFSR[7] ^~ LFSR[6];
            // end
            // 8: begin
            //     r_XNOR = LFSR[8] ^~ LFSR[6] ^~ LFSR[5] ^~ LFSR[4];
            // end
            // 9: begin
            //     r_XNOR = LFSR[9] ^~ LFSR[5];
            // end
            // 10: begin
            //     r_XNOR = LFSR[10] ^~ LFSR[7];
            // end
            // 11: begin
            //     r_XNOR = LFSR[11] ^~ LFSR[9];
            // end
            // 12: begin
            //     r_XNOR = LFSR[12] ^~ LFSR[6] ^~ LFSR[4] ^~ LFSR[1];
            // end
            // 13: begin
            //     r_XNOR = LFSR[13] ^~ LFSR[4] ^~ LFSR[3] ^~ LFSR[1];
            // end
            // 14: begin
            //     r_XNOR = LFSR[14] ^~ LFSR[5] ^~ LFSR[3] ^~ LFSR[1];
            // end
            // 15: begin
            //     r_XNOR = LFSR[15] ^~ LFSR[14];
            // end
            // 16: begin
            //     r_XNOR = LFSR[16] ^~ LFSR[15] ^~ LFSR[13] ^~ LFSR[4];
            // end
            // 17: begin
            //     r_XNOR = LFSR[17] ^~ LFSR[14];
            // end
            // 18: begin
            //     r_XNOR = LFSR[18] ^~ LFSR[11];
            // end
            // 19: begin
            //     r_XNOR = LFSR[19] ^~ LFSR[6] ^~ LFSR[2] ^~ LFSR[1];
            // end
            // 20: begin
            //     r_XNOR = LFSR[20] ^~ LFSR[17];
            // end
            // 21: begin
            //     r_XNOR = LFSR[21] ^~ LFSR[19];
            // end
            // 22: begin
            //     r_XNOR = LFSR[22] ^~ LFSR[21];
            // end
            // 23: begin
            //     r_XNOR = LFSR[23] ^~ LFSR[18];
            // end
            // 24: begin
            //     r_XNOR = LFSR[24] ^~ LFSR[23] ^~ LFSR[22] ^~ LFSR[17];
            // end
            // 25: begin
            //     r_XNOR = LFSR[25] ^~ LFSR[22];
            // end
            // 26: begin
            //     r_XNOR = LFSR[26] ^~ LFSR[6] ^~ LFSR[2] ^~ LFSR[1];
            // end
            // 27: begin
            //     r_XNOR = LFSR[27] ^~ LFSR[5] ^~ LFSR[2] ^~ LFSR[1];
            // end
            // 28: begin
            //     r_XNOR = LFSR[28] ^~ LFSR[25];
            // end
            // 29: begin
            //     r_XNOR = LFSR[29] ^~ LFSR[27];
            // end
            // 30: begin
            //     r_XNOR = LFSR[30] ^~ LFSR[6] ^~ LFSR[4] ^~ LFSR[1];
            // end
            // 31: begin
            //     r_XNOR = LFSR[31] ^~ LFSR[28];
            // end
            // 32: begin
            //     r_XNOR = LFSR[32] ^~ LFSR[22] ^~ LFSR[2] ^~ LFSR[1];
            // end
        endcase
    end

    assign data_out = LFSR;

endmodule

