`include "sys_defs.svh"

module stage_issue (
    input clock,
    input reset,
    input logic mispredict,

    input RS_BANKS rs_banks,                                  // Structured RS entries
    input FU_GRANTS fu_grants,                                // FU availability (structured)

    output ISSUE_CLEAR issue_clear,                           // Clear signals (structured)
    output ISSUE_ENTRIES issue_entries                        // To EX stage (structured)
);

    // Helper: Check if RS entry is ready
    function automatic logic is_ready(RS_ENTRY entry);
        return entry.valid && entry.src1_ready && entry.src2_ready;
    endfunction

    // Internal state (structured)
    ISSUE_ENTRIES issue_register, issue_register_next;

    // Ready signals for each RS bank
    logic [`RS_ALU_SZ-1:0]    rs_ready_alu;
    logic [`RS_MULT_SZ-1:0]   rs_ready_mult;
    logic [`RS_BRANCH_SZ-1:0] rs_ready_branch;
    logic [`RS_MEM_SZ-1:0]    rs_ready_mem;

    // Grant outputs from allocators
    logic [`NUM_FU_ALU-1:0][`RS_ALU_SZ-1:0] grants_alu;
    logic [`NUM_FU_MULT-1:0][`RS_MULT_SZ-1:0] grants_mult;
    logic [`NUM_FU_BRANCH-1:0][`RS_BRANCH_SZ-1:0] grants_branch;
    logic [`NUM_FU_MEM-1:0][`RS_MEM_SZ-1:0] grants_mem;

    // Compute ready signals for each bank
    always_comb begin
        for (int i = 0; i < `RS_ALU_SZ; i++) begin
            rs_ready_alu[i] = is_ready(rs_banks.alu[i]);
        end
        for (int i = 0; i < `RS_MULT_SZ; i++) begin
            rs_ready_mult[i] = is_ready(rs_banks.mult[i]);
        end
        for (int i = 0; i < `RS_BRANCH_SZ; i++) begin
            rs_ready_branch[i] = is_ready(rs_banks.branch[i]);
        end
        for (int i = 0; i < `RS_MEM_SZ; i++) begin
            rs_ready_mem[i] = is_ready(rs_banks.mem[i]);
        end
    end

    // Allocators for each FU category
    allocator #(.NUM_RESOURCES(`RS_ALU_SZ), .NUM_REQUESTS(`NUM_FU_ALU)) alu_allocator (
        .reset(reset | mispredict), .clock(clock),
        .req(rs_ready_alu),
        .clear(fu_grants.alu),
        .grant(grants_alu)
    );

    allocator #(.NUM_RESOURCES(`RS_MULT_SZ), .NUM_REQUESTS(`NUM_FU_MULT)) mult_allocator (
        .reset(reset | mispredict), .clock(clock),
        .req(rs_ready_mult),
        .clear(fu_grants.mult),
        .grant(grants_mult)
    );

    allocator #(.NUM_RESOURCES(`RS_BRANCH_SZ), .NUM_REQUESTS(`NUM_FU_BRANCH)) branch_allocator (
        .reset(reset | mispredict), .clock(clock),
        .req(rs_ready_branch),
        .clear(fu_grants.branch),
        .grant(grants_branch)
    );

    allocator #(.NUM_RESOURCES(`RS_MEM_SZ), .NUM_REQUESTS(`NUM_FU_MEM)) mem_allocator (
        .reset(reset | mispredict), .clock(clock),
        .req(rs_ready_mem),
        .clear(fu_grants.mem),
        .grant(grants_mem)
    );

    // Generate clear signals (grant to index conversion)
    // Note: clear indices contain local RS bank indices since each RS module
    // maintains its own entry array. The RS modules handle their own indexing.
    always_comb begin
        issue_clear = '0;

        // ALU - use local ALU RS indices
        for (int fu = 0; fu < `NUM_FU_ALU; fu++) begin
            for (int rs = 0; rs < `RS_ALU_SZ; rs++) begin
                if (grants_alu[fu][rs]) begin
                    issue_clear.valid_alu[fu] = 1'b1;
                    issue_clear.idxs_alu[fu] = RS_IDX'(rs);
                end
            end
        end

        // MULT - use local MULT RS indices
        for (int fu = 0; fu < `NUM_FU_MULT; fu++) begin
            for (int rs = 0; rs < `RS_MULT_SZ; rs++) begin
                if (grants_mult[fu][rs]) begin
                    issue_clear.valid_mult[fu] = 1'b1;
                    issue_clear.idxs_mult[fu] = RS_IDX'(rs);
                end
            end
        end

        // BRANCH - use local BRANCH RS indices
        for (int fu = 0; fu < `NUM_FU_BRANCH; fu++) begin
            for (int rs = 0; rs < `RS_BRANCH_SZ; rs++) begin
                if (grants_branch[fu][rs]) begin
                    issue_clear.valid_branch[fu] = 1'b1;
                    issue_clear.idxs_branch[fu] = RS_IDX'(rs);
                end
            end
        end

        // MEM - use local MEM RS indices
        for (int fu = 0; fu < `NUM_FU_MEM; fu++) begin
            for (int rs = 0; rs < `RS_MEM_SZ; rs++) begin
                if (grants_mem[fu][rs]) begin
                    issue_clear.valid_mem[fu] = 1'b1;
                    issue_clear.idxs_mem[fu] = RS_IDX'(rs);
                end
            end
        end
    end

    // Update issue register from granted RS entries
    always_comb begin
        issue_register_next = issue_register;

        // ALU - use structured ALU bank
        for (int fu = 0; fu < `NUM_FU_ALU; fu++) begin
            if (fu_grants.alu[fu]) begin
                for (int rs = 0; rs < `RS_ALU_SZ; rs++) begin
                    if (grants_alu[fu][rs]) begin
                        issue_register_next.alu[fu] = rs_banks.alu[rs];
                    end
                end
            end
        end

        // MULT - use structured MULT bank
        for (int fu = 0; fu < `NUM_FU_MULT; fu++) begin
            if (fu_grants.mult[fu]) begin
                for (int rs = 0; rs < `RS_MULT_SZ; rs++) begin
                    if (grants_mult[fu][rs]) begin
                        issue_register_next.mult[fu] = rs_banks.mult[rs];
                    end
                end
            end
        end

        // BRANCH - use structured BRANCH bank
        for (int fu = 0; fu < `NUM_FU_BRANCH; fu++) begin
            if (fu_grants.branch[fu]) begin
                for (int rs = 0; rs < `RS_BRANCH_SZ; rs++) begin
                    if (grants_branch[fu][rs]) begin
                        issue_register_next.branch[fu] = rs_banks.branch[rs];
                    end
                end
            end
        end

        // MEM - use structured MEM bank
        for (int fu = 0; fu < `NUM_FU_MEM; fu++) begin
            if (fu_grants.mem[fu]) begin
                for (int rs = 0; rs < `RS_MEM_SZ; rs++) begin
                    if (grants_mem[fu][rs]) begin
                        issue_register_next.mem[fu] = rs_banks.mem[rs];
                    end
                end
            end
        end
    end

    // Output assignment
    assign issue_entries = issue_register;

    always_ff @(posedge clock) begin
        if (reset | mispredict) begin
            issue_register <= '0;
        end else begin
            issue_register <= issue_register_next;
        end
    end

endmodule
